`default_nettype none

module uart #(
    parameter DELAY_FRAMES = 234  // 27,000,000 (27Mhz) / 115200 Baud rate
) (
    input clk,
    input uartRx,
    output reg byteReady,
    output reg [7:0] dataIn
);

  localparam HALF_DELAY_WAIT = (DELAY_FRAMES / 2);

  reg [ 3:0] rxState = 0;
  reg [12:0] rxCounter = 0;
  reg [ 2:0] rxBitNumber = 0;

  localparam RX_STATE_IDLE = 0;
  localparam RX_STATE_START_BIT = 1;
  localparam RX_STATE_READ_WAIT = 2;
  localparam RX_STATE_READ = 3;
  localparam RX_STATE_STOP_BIT = 5;

  always @(posedge clk) begin
    case (rxState)
      RX_STATE_IDLE: begin
        if (uartRx == 0) begin
          rxState <= RX_STATE_START_BIT;
          rxCounter <= 1;
          rxBitNumber <= 0;
          byteReady <= 0;
        end
      end
      RX_STATE_START_BIT: begin
        if (rxCounter == HALF_DELAY_WAIT) begin
          rxState   <= RX_STATE_READ_WAIT;
          rxCounter <= 1;
        end else rxCounter <= rxCounter + 1;
      end
      RX_STATE_READ_WAIT: begin
        rxCounter <= rxCounter + 1;
        if ((rxCounter + 1) == DELAY_FRAMES) begin
          rxState <= RX_STATE_READ;
        end
      end
      RX_STATE_READ: begin
        rxCounter <= 1;
        dataIn <= {uartRx, dataIn[7:1]};
        rxBitNumber <= rxBitNumber + 1;
        if (rxBitNumber == 3'b111) rxState <= RX_STATE_STOP_BIT;
        else rxState <= RX_STATE_READ_WAIT;
      end
      RX_STATE_STOP_BIT: begin
        rxCounter <= rxCounter + 1;
        if ((rxCounter + 1) == DELAY_FRAMES) begin
          rxState   <= RX_STATE_IDLE;
          rxCounter <= 0;
          byteReady <= 1;
        end
      end
    endcase
  end
endmodule
